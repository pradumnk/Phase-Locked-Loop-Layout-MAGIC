magic
tech scmos
timestamp 1647145390
<< nwell >>
rect -1148 69 -1116 112
rect -103 65 -71 108
rect -41 65 -9 108
rect 13 65 45 108
rect 76 65 108 108
rect -1381 -16 -1349 27
rect -1290 -16 -1258 27
rect -41 20 -9 52
rect 14 20 46 52
rect 76 21 108 53
rect -1148 -147 -1116 -104
rect -413 -115 -346 -80
<< polysilicon >>
rect -1135 121 -1083 127
rect -1397 96 -1195 102
rect -1135 98 -1131 121
rect -1397 9 -1392 96
rect -1135 77 -1131 82
rect -1135 60 -1131 65
rect -1397 3 -1371 9
rect -1360 3 -1356 9
rect -1397 -22 -1392 3
rect -1311 0 -1280 7
rect -1269 0 -1263 7
rect -1397 -122 -1392 -33
rect -1397 -129 -1371 -122
rect -1360 -129 -1356 -122
rect -1311 -125 -1306 0
rect -1135 -52 -1131 44
rect -1200 -59 -1131 -52
rect -1135 -119 -1131 -59
rect -1311 -132 -1280 -125
rect -1269 -132 -1264 -125
rect -1311 -183 -1306 -132
rect -1135 -138 -1131 -135
rect -1087 -164 -1083 121
rect -92 88 94 92
rect -92 84 -86 88
rect -28 83 -22 88
rect -92 45 -86 72
rect 27 82 33 88
rect 88 82 94 88
rect -28 66 -22 71
rect 27 65 33 70
rect 88 65 94 70
rect -30 43 -23 47
rect 27 43 34 47
rect 88 43 95 47
rect -30 3 -23 31
rect 27 7 34 31
rect 88 7 95 31
rect -126 -7 -23 3
rect 11 -2 34 7
rect 71 -2 95 7
rect -30 -13 -23 -7
rect 27 -13 34 -2
rect 88 -13 95 -2
rect -30 -30 -23 -25
rect 27 -30 34 -25
rect 88 -30 95 -25
rect -687 -65 -603 -40
rect -687 -90 -678 -65
rect -91 -70 -85 -64
rect -29 -70 -23 -63
rect 28 -69 34 -63
rect 89 -69 95 -63
rect -391 -90 -382 -83
rect -91 -86 -85 -82
rect -29 -86 -23 -82
rect 0 -86 7 -85
rect 28 -86 34 -81
rect 89 -86 95 -81
rect -687 -95 -582 -90
rect -590 -105 -582 -95
rect -687 -109 -582 -105
rect -91 -92 95 -86
rect -687 -119 -678 -109
rect -687 -125 -582 -119
rect -391 -120 -382 -107
rect -591 -144 -582 -125
rect -398 -131 -382 -120
rect 0 -127 7 -92
rect -391 -137 -382 -131
rect -685 -149 -582 -144
rect -685 -159 -678 -149
rect -685 -163 -582 -159
rect -391 -161 -382 -154
rect -588 -173 -582 -163
rect -1087 -183 -1083 -176
rect -1311 -188 -1083 -183
rect -685 -181 -582 -173
rect -685 -199 -673 -181
rect -685 -223 -599 -199
<< ndiffusion >>
rect -1145 56 -1135 60
rect -1145 48 -1143 56
rect -1137 48 -1135 56
rect -1145 44 -1135 48
rect -1131 56 -1119 60
rect -1131 48 -1128 56
rect -1122 48 -1119 56
rect -1131 44 -1119 48
rect -1371 -110 -1360 -109
rect -1371 -116 -1368 -110
rect -1363 -116 -1360 -110
rect -1371 -122 -1360 -116
rect -1280 -113 -1269 -112
rect -1280 -119 -1277 -113
rect -1272 -119 -1269 -113
rect -1280 -125 -1269 -119
rect -1371 -135 -1360 -129
rect -1371 -141 -1368 -135
rect -1363 -141 -1360 -135
rect -1280 -137 -1269 -132
rect -1280 -143 -1277 -137
rect -1272 -143 -1269 -137
rect -1280 -144 -1269 -143
rect -1145 -161 -1119 -157
rect -1145 -169 -1143 -161
rect -1137 -169 -1128 -161
rect -1122 -169 -1119 -161
rect -1145 -173 -1119 -169
rect -37 -16 -30 -13
rect -37 -23 -36 -16
rect -32 -23 -30 -16
rect -37 -25 -30 -23
rect -23 -16 -15 -13
rect -23 -23 -20 -16
rect -16 -23 -15 -16
rect -23 -25 -15 -23
rect 19 -16 27 -13
rect 19 -23 20 -16
rect 24 -23 27 -16
rect 19 -25 27 -23
rect 34 -16 41 -13
rect 34 -23 36 -16
rect 40 -23 41 -16
rect 34 -25 41 -23
rect 81 -16 88 -13
rect 81 -23 82 -16
rect 86 -23 88 -16
rect 81 -25 88 -23
rect 95 -16 103 -13
rect 95 -23 98 -16
rect 102 -23 103 -16
rect 95 -25 103 -23
rect -98 -73 -91 -70
rect -98 -80 -97 -73
rect -93 -80 -91 -73
rect -98 -82 -91 -80
rect -85 -73 -76 -70
rect -85 -80 -82 -73
rect -78 -80 -76 -73
rect -85 -82 -76 -80
rect -37 -73 -29 -70
rect -37 -80 -35 -73
rect -31 -80 -29 -73
rect -37 -82 -29 -80
rect -23 -73 -15 -70
rect -23 -80 -21 -73
rect -17 -80 -15 -73
rect -23 -82 -15 -80
rect 20 -72 28 -69
rect 20 -79 21 -72
rect 25 -79 28 -72
rect 20 -81 28 -79
rect 34 -72 42 -69
rect 34 -79 37 -72
rect 41 -79 42 -72
rect 34 -81 42 -79
rect 81 -72 89 -69
rect 81 -79 82 -72
rect 86 -79 89 -72
rect 81 -81 89 -79
rect 95 -72 103 -69
rect 95 -79 98 -72
rect 102 -79 103 -72
rect 95 -81 103 -79
rect -403 -154 -391 -137
rect -382 -139 -356 -137
rect -382 -151 -372 -139
rect -363 -151 -356 -139
rect -382 -154 -356 -151
<< pdiffusion >>
rect -1145 93 -1135 98
rect -1145 85 -1143 93
rect -1137 85 -1135 93
rect -1145 82 -1135 85
rect -1131 93 -1119 98
rect -1131 85 -1128 93
rect -1122 85 -1119 93
rect -1131 82 -1119 85
rect -1371 20 -1360 21
rect -1371 13 -1368 20
rect -1363 13 -1360 20
rect -1371 9 -1360 13
rect -1280 19 -1269 21
rect -1280 12 -1277 19
rect -1272 12 -1269 19
rect -1280 7 -1269 12
rect -1371 -3 -1360 3
rect -1371 -10 -1368 -3
rect -1363 -10 -1360 -3
rect -1371 -11 -1360 -10
rect -1280 -4 -1269 0
rect -1280 -11 -1277 -4
rect -1272 -11 -1269 -4
rect -1145 -125 -1135 -119
rect -1145 -133 -1143 -125
rect -1137 -133 -1135 -125
rect -1145 -135 -1135 -133
rect -1131 -125 -1119 -119
rect -1131 -133 -1128 -125
rect -1122 -133 -1119 -125
rect -1131 -135 -1119 -133
rect -98 82 -92 84
rect -98 74 -97 82
rect -93 74 -92 82
rect -98 72 -92 74
rect -86 82 -76 84
rect -86 75 -82 82
rect -78 75 -76 82
rect -86 72 -76 75
rect -37 80 -28 83
rect -37 73 -36 80
rect -31 73 -28 80
rect -37 71 -28 73
rect -22 81 -15 83
rect -22 73 -21 81
rect -16 73 -15 81
rect -22 71 -15 73
rect 18 79 27 82
rect 18 72 20 79
rect 24 72 27 79
rect 18 70 27 72
rect 33 79 40 82
rect 33 72 35 79
rect 39 72 40 79
rect 33 70 40 72
rect 81 79 88 82
rect 81 72 82 79
rect 87 72 88 79
rect 81 70 88 72
rect 94 79 103 82
rect 94 72 97 79
rect 101 72 103 79
rect 94 70 103 72
rect -37 40 -30 43
rect -37 33 -36 40
rect -32 33 -30 40
rect -37 31 -30 33
rect -23 40 -15 43
rect -23 33 -20 40
rect -16 33 -15 40
rect -23 31 -15 33
rect 19 40 27 43
rect 19 33 20 40
rect 24 33 27 40
rect 19 31 27 33
rect 34 40 41 43
rect 34 33 36 40
rect 40 33 41 40
rect 34 31 41 33
rect 81 40 88 43
rect 81 33 82 40
rect 86 33 88 40
rect 81 31 88 33
rect 95 40 103 43
rect 95 33 97 40
rect 102 33 103 40
rect 95 31 103 33
rect -403 -107 -391 -90
rect -382 -94 -356 -90
rect -382 -106 -372 -94
rect -363 -106 -356 -94
rect -382 -107 -356 -106
<< metal1 >>
rect 140 212 159 213
rect -159 206 159 212
rect -1057 188 159 206
rect -1195 71 -1189 96
rect -1143 71 -1137 85
rect -1195 63 -1137 71
rect -1368 59 -1272 60
rect -1368 53 -1361 59
rect -1356 53 -1337 59
rect -1332 53 -1294 59
rect -1289 53 -1272 59
rect -1368 52 -1272 53
rect -1368 20 -1363 52
rect -1277 19 -1272 52
rect -1143 56 -1137 63
rect -1128 56 -1122 85
rect -1449 -33 -1398 -22
rect -1368 -58 -1363 -10
rect -1422 -71 -1363 -58
rect -1422 -199 -1413 -71
rect -1368 -110 -1363 -71
rect -1277 -49 -1272 -11
rect -1277 -52 -1195 -49
rect -1277 -59 -1206 -52
rect -1200 -59 -1195 -52
rect -1277 -62 -1195 -59
rect -1277 -113 -1272 -62
rect -1128 -125 -1122 48
rect -1368 -163 -1363 -141
rect -1277 -163 -1272 -143
rect -1368 -168 -1358 -163
rect -1354 -168 -1340 -163
rect -1336 -168 -1296 -163
rect -1292 -168 -1272 -163
rect -1143 -161 -1137 -133
rect -1143 -199 -1137 -169
rect -1422 -210 -1137 -199
rect -1128 -161 -1122 -133
rect -1057 -164 -1050 188
rect -159 187 159 188
rect -159 9 -141 187
rect -100 103 105 104
rect -100 102 -38 103
rect -96 97 -90 102
rect -86 97 -81 102
rect -77 98 -38 102
rect -34 98 -30 103
rect -26 98 -15 103
rect -11 98 15 103
rect 19 98 24 103
rect 28 98 40 103
rect 44 98 78 103
rect 82 98 87 103
rect 91 98 100 103
rect 104 98 105 103
rect -77 97 105 98
rect -97 82 -93 97
rect -21 81 -16 97
rect -82 45 -78 75
rect -159 3 -126 9
rect -772 -22 -583 3
rect -159 -7 -132 3
rect -159 -14 -126 -7
rect -1128 -208 -1122 -169
rect -1083 -176 -1050 -164
rect -770 -208 -757 -22
rect -603 -40 -584 -22
rect -82 -73 -78 39
rect 35 79 39 97
rect 97 79 100 97
rect -36 40 -32 73
rect 20 40 24 72
rect 82 40 86 72
rect -20 9 -16 33
rect 36 9 40 33
rect -20 7 11 9
rect -20 -2 5 7
rect -20 -4 11 -2
rect 36 7 71 9
rect 36 -2 65 7
rect 36 -4 71 -2
rect 98 8 102 33
rect 140 8 159 187
rect 98 -3 180 8
rect -20 -16 -16 -4
rect 36 -16 40 -4
rect 98 -16 102 -3
rect -35 -73 -32 -23
rect 21 -72 24 -23
rect 82 -72 86 -23
rect -372 -120 -363 -106
rect -97 -104 -93 -80
rect -21 -104 -17 -80
rect 37 -104 41 -79
rect -97 -111 -91 -104
rect -86 -111 -77 -104
rect -72 -111 -64 -104
rect -59 -111 -38 -104
rect -33 -111 -26 -104
rect -21 -111 -10 -104
rect -5 -111 14 -104
rect 19 -111 28 -104
rect 33 -111 46 -104
rect 51 -111 59 -104
rect 64 -111 73 -104
rect 78 -111 93 -104
rect 98 -111 102 -79
rect -509 -131 -405 -120
rect -372 -131 -371 -120
rect -364 -131 -363 -120
rect -509 -132 -419 -131
rect -508 -199 -496 -132
rect -372 -139 -363 -131
rect -372 -152 -363 -151
rect -1128 -221 -757 -208
rect -1128 -222 -758 -221
rect -582 -200 -496 -199
rect 0 -200 7 -139
rect -582 -223 7 -200
rect -507 -224 7 -223
<< ntransistor >>
rect -1135 44 -1131 60
rect -1371 -129 -1360 -122
rect -1280 -132 -1269 -125
rect -30 -25 -23 -13
rect 27 -25 34 -13
rect 88 -25 95 -13
rect -91 -82 -85 -70
rect -29 -82 -23 -70
rect 28 -81 34 -69
rect 89 -81 95 -69
rect -391 -154 -382 -137
<< ptransistor >>
rect -1135 82 -1131 98
rect -1371 3 -1360 9
rect -1280 0 -1269 7
rect -1135 -135 -1131 -119
rect -92 72 -86 84
rect -28 71 -22 83
rect 27 70 33 82
rect 88 70 94 82
rect -30 31 -23 43
rect 27 31 34 43
rect 88 31 95 43
rect -391 -107 -382 -90
<< polycontact >>
rect -1195 96 -1189 102
rect -1398 -33 -1392 -22
rect -1206 -59 -1200 -52
rect -92 39 -78 45
rect -132 -7 -126 3
rect 5 -2 11 7
rect 65 -2 71 7
rect -603 -65 -584 -40
rect -405 -131 -398 -120
rect 0 -139 7 -127
rect -1087 -176 -1083 -164
rect -599 -223 -582 -199
<< ndcontact >>
rect -1143 48 -1137 56
rect -1128 48 -1122 56
rect -1368 -116 -1363 -110
rect -1277 -119 -1272 -113
rect -1368 -141 -1363 -135
rect -1277 -143 -1272 -137
rect -1143 -169 -1137 -161
rect -1128 -169 -1122 -161
rect -36 -23 -32 -16
rect -20 -23 -16 -16
rect 20 -23 24 -16
rect 36 -23 40 -16
rect 82 -23 86 -16
rect 98 -23 102 -16
rect -97 -80 -93 -73
rect -82 -80 -78 -73
rect -35 -80 -31 -73
rect -21 -80 -17 -73
rect 21 -79 25 -72
rect 37 -79 41 -72
rect 82 -79 86 -72
rect 98 -79 102 -72
rect -372 -151 -363 -139
<< pdcontact >>
rect -1143 85 -1137 93
rect -1128 85 -1122 93
rect -1368 13 -1363 20
rect -1277 12 -1272 19
rect -1368 -10 -1363 -3
rect -1277 -11 -1272 -4
rect -1143 -133 -1137 -125
rect -1128 -133 -1122 -125
rect -97 74 -93 82
rect -82 75 -78 82
rect -36 73 -31 80
rect -21 73 -16 81
rect 20 72 24 79
rect 35 72 39 79
rect 82 72 87 79
rect 97 72 101 79
rect -36 33 -32 40
rect -20 33 -16 40
rect 20 33 24 40
rect 36 33 40 40
rect 82 33 86 40
rect 97 33 102 40
rect -372 -106 -363 -94
<< psubstratepcontact >>
rect -1358 -168 -1354 -163
rect -1340 -168 -1336 -163
rect -1296 -168 -1292 -163
rect -91 -111 -86 -104
rect -77 -111 -72 -104
rect -64 -111 -59 -104
rect -38 -111 -33 -104
rect -26 -111 -21 -104
rect -10 -111 -5 -104
rect -371 -131 -364 -120
rect 14 -111 19 -104
rect 28 -111 33 -104
rect 46 -111 51 -104
rect 59 -111 64 -104
rect 73 -111 78 -104
rect 93 -111 98 -104
<< nsubstratencontact >>
rect -1361 53 -1356 59
rect -1337 53 -1332 59
rect -1294 53 -1289 59
rect -100 97 -96 102
rect -90 97 -86 102
rect -81 97 -77 102
rect -38 98 -34 103
rect -30 98 -26 103
rect -15 98 -11 103
rect 15 98 19 103
rect 24 98 28 103
rect 40 98 44 103
rect 78 98 82 103
rect 87 98 91 103
rect 100 98 104 103
<< labels >>
rlabel metal1 -100 103 -99 103 5 vdd
rlabel metal1 2 -155 3 -155 1 vctrl
rlabel metal1 128 1 129 1 1 out
rlabel metal1 -96 -109 -96 -109 1 gnd
rlabel metal1 -82 7 -82 7 1 mid1
rlabel metal1 -11 2 -11 2 1 mid2
rlabel metal1 43 1 43 1 1 mid3
rlabel metal1 -35 58 -35 58 1 top1
rlabel metal1 21 58 21 58 1 top2
rlabel metal1 83 58 83 58 1 top3
rlabel metal1 -34 -50 -34 -50 1 bot1
rlabel metal1 21 -47 21 -47 1 bot2
rlabel metal1 83 -48 83 -48 1 bot3
rlabel metal1 -1367 58 -1367 58 1 vdd
rlabel metal1 -1367 -165 -1367 -165 1 gnd
rlabel metal1 -371 -133 -371 -133 1 gnd
rlabel metal1 -1446 -28 -1446 -28 3 ip
rlabel metal1 -1367 -54 -1367 -54 1 ip_bar
rlabel metal1 -1276 -50 -1276 -50 1 ip2_bar
rlabel metal1 -1037 -219 -1037 -219 1 op_xor
rlabel metal1 -1192 66 -1192 66 1 net1
<< end >>
