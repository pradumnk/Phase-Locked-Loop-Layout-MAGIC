* SPICE3 file created from vco.ext - technology: scmos

.include model_VlsiDesign.txt 

.param Lmin=0.4U
.param Wn=1.009U
.param Wp=2.435U

M1000 mid1 mid1 vdd vdd cmosp        L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1001 mid2 out bot1 gnd cmosn        L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1002 vdd mid1 top1 vdd cmosp        L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1003 mid1 vctrl gnd gnd cmosn       L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1004 gnd vctrl bot1 gnd cmosn       L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1005 out mid3 top3 w_76_21 cmosp   L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1006 out mid3 bot3 gnd cmosn        L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1007 vdd mid1 top3 vdd cmosp        L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1008 mid3 mid2 bot2 gnd cmosn       L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1009 gnd vctrl bot3 gnd cmosn       L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1010 gnd vctrl bot2 gnd cmosn       L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1011 mid2 out top1 w_n41_20 cmosp  L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1012 mid3 mid2 top2 w_14_20 cmosp  L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1013 vdd mid1 top2 vdd cmosp        L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1014 net1 ip vdd vdd cmosp          L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1015 net1 ip gnd gnd cmosn          L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1016 out_xor out ip ip cmosp        L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1017 out_xor out net1 net1 cmosn    L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
M1018 out ip out_xor out_xor cmosp   L=Lmin W=Wp AD=(2*Lmin*Wp) AS=(2*Lmin*Wp) PD=(2*Wp+4*Lmin) PS=(2*Wp+4*Lmin)
M1019 out net1 out_xor out_xor cmosn L=Lmin W=Wn AD =(2*wn*lmin) AS =(2*wn*lmin) PD =(2*wn+4*lmin) PS =(2*wn+4*lmin)
C0 mid3 w_14_20 2.07fF
C1 mid2 w_14_20 8.18fF
C2 mid1 vdd 54.93fF
C3 vctrl gnd 2.91fF
C4 w_n41_20 out 8.18fF
C5 w_76_21 mid3 7.74fF
C6 w_n41_20 mid2 2.07fF
R19 out_xor vctrl 0.00000000005
C7 gnd gnd 58.09fF
C8 vctrl gnd 102.72fF
C9 bot3 gnd 8.27fF
C10 bot2 gnd 6.20fF
C11 bot1 gnd 6.34fF
C12 mid3 gnd 52.93fF
C13 mid2 gnd 49.54fF
C14 out gnd 1.11fF
C15 top2 gnd 2.44fF
C16 top1 gnd 2.44fF
C17 mid1 gnd 100.44fF
C18 vdd gnd 7.31fF
v1 vdd gnd 3.3
vip ip gnd dc 0 pulse(0 3.3 4ns 2ps 2ps 1.8ns 3ns)

.tran 1ns 150ns 0ns
.control
run
plot v(ip) v(out)
.endc
.end