magic
tech scmos
timestamp 1646889068
<< nwell >>
rect -103 65 -71 108
rect -41 65 -9 108
rect 13 65 45 108
rect 76 65 108 108
rect -41 20 -9 52
rect 14 20 46 52
rect 76 21 108 53
<< polysilicon >>
rect -92 88 94 92
rect -92 84 -86 88
rect -28 83 -22 88
rect -92 45 -86 72
rect 27 82 33 88
rect 88 82 94 88
rect -28 66 -22 71
rect 27 65 33 70
rect 88 65 94 70
rect -30 43 -23 47
rect 27 43 34 47
rect 88 43 95 47
rect -30 3 -23 31
rect 27 7 34 31
rect 88 7 95 31
rect -126 -7 -23 3
rect 11 -2 34 7
rect 71 -2 95 7
rect -30 -13 -23 -7
rect 27 -13 34 -2
rect 88 -13 95 -2
rect -30 -30 -23 -25
rect 27 -30 34 -25
rect 88 -30 95 -25
rect -91 -70 -85 -64
rect -29 -70 -23 -63
rect 28 -69 34 -63
rect 89 -69 95 -63
rect -91 -86 -85 -82
rect -29 -86 -23 -82
rect 0 -86 7 -85
rect 28 -86 34 -81
rect 89 -86 95 -81
rect -91 -92 95 -86
rect 0 -127 7 -92
<< ndiffusion >>
rect -37 -16 -30 -13
rect -37 -23 -36 -16
rect -32 -23 -30 -16
rect -37 -25 -30 -23
rect -23 -16 -15 -13
rect -23 -23 -20 -16
rect -16 -23 -15 -16
rect -23 -25 -15 -23
rect 19 -16 27 -13
rect 19 -23 20 -16
rect 24 -23 27 -16
rect 19 -25 27 -23
rect 34 -16 41 -13
rect 34 -23 36 -16
rect 40 -23 41 -16
rect 34 -25 41 -23
rect 81 -16 88 -13
rect 81 -23 82 -16
rect 86 -23 88 -16
rect 81 -25 88 -23
rect 95 -16 103 -13
rect 95 -23 98 -16
rect 102 -23 103 -16
rect 95 -25 103 -23
rect -98 -73 -91 -70
rect -98 -80 -97 -73
rect -93 -80 -91 -73
rect -98 -82 -91 -80
rect -85 -73 -76 -70
rect -85 -80 -82 -73
rect -78 -80 -76 -73
rect -85 -82 -76 -80
rect -37 -73 -29 -70
rect -37 -80 -35 -73
rect -31 -80 -29 -73
rect -37 -82 -29 -80
rect -23 -73 -15 -70
rect -23 -80 -21 -73
rect -17 -80 -15 -73
rect -23 -82 -15 -80
rect 20 -72 28 -69
rect 20 -79 21 -72
rect 25 -79 28 -72
rect 20 -81 28 -79
rect 34 -72 42 -69
rect 34 -79 37 -72
rect 41 -79 42 -72
rect 34 -81 42 -79
rect 81 -72 89 -69
rect 81 -79 82 -72
rect 86 -79 89 -72
rect 81 -81 89 -79
rect 95 -72 103 -69
rect 95 -79 98 -72
rect 102 -79 103 -72
rect 95 -81 103 -79
<< pdiffusion >>
rect -98 82 -92 84
rect -98 74 -97 82
rect -93 74 -92 82
rect -98 72 -92 74
rect -86 82 -76 84
rect -86 75 -82 82
rect -78 75 -76 82
rect -86 72 -76 75
rect -37 80 -28 83
rect -37 73 -36 80
rect -31 73 -28 80
rect -37 71 -28 73
rect -22 81 -15 83
rect -22 73 -21 81
rect -16 73 -15 81
rect -22 71 -15 73
rect 18 79 27 82
rect 18 72 20 79
rect 24 72 27 79
rect 18 70 27 72
rect 33 79 40 82
rect 33 72 35 79
rect 39 72 40 79
rect 33 70 40 72
rect 81 79 88 82
rect 81 72 82 79
rect 87 72 88 79
rect 81 70 88 72
rect 94 79 103 82
rect 94 72 97 79
rect 101 72 103 79
rect 94 70 103 72
rect -37 40 -30 43
rect -37 33 -36 40
rect -32 33 -30 40
rect -37 31 -30 33
rect -23 40 -15 43
rect -23 33 -20 40
rect -16 33 -15 40
rect -23 31 -15 33
rect 19 40 27 43
rect 19 33 20 40
rect 24 33 27 40
rect 19 31 27 33
rect 34 40 41 43
rect 34 33 36 40
rect 40 33 41 40
rect 34 31 41 33
rect 81 40 88 43
rect 81 33 82 40
rect 86 33 88 40
rect 81 31 88 33
rect 95 40 103 43
rect 95 33 97 40
rect 102 33 103 40
rect 95 31 103 33
<< metal1 >>
rect -100 103 105 104
rect -100 102 -38 103
rect -96 97 -90 102
rect -86 97 -81 102
rect -77 98 -38 102
rect -34 98 -30 103
rect -26 98 -15 103
rect -11 98 15 103
rect 19 98 24 103
rect 28 98 40 103
rect 44 98 78 103
rect 82 98 87 103
rect 91 98 100 103
rect 104 98 105 103
rect -77 97 105 98
rect -97 82 -93 97
rect -21 81 -16 97
rect -82 45 -78 75
rect -159 3 -126 9
rect -159 -7 -132 3
rect -159 -14 -126 -7
rect -159 -188 -143 -14
rect -82 -73 -78 39
rect 35 79 39 97
rect 97 79 100 97
rect -36 40 -32 73
rect 20 40 24 72
rect 82 40 86 72
rect -20 9 -16 33
rect 36 9 40 33
rect -20 7 11 9
rect -20 -2 5 7
rect -20 -4 11 -2
rect 36 7 71 9
rect 36 -2 65 7
rect 36 -4 71 -2
rect 98 8 102 33
rect 98 -3 180 8
rect -20 -16 -16 -4
rect 36 -16 40 -4
rect 98 -16 102 -3
rect -35 -73 -32 -23
rect 21 -72 24 -23
rect 82 -72 86 -23
rect -97 -104 -93 -80
rect -21 -104 -17 -80
rect 37 -104 41 -79
rect -97 -111 -91 -104
rect -86 -111 -77 -104
rect -72 -111 -64 -104
rect -59 -111 -38 -104
rect -33 -111 -26 -104
rect -21 -111 -10 -104
rect -5 -111 14 -104
rect 19 -111 28 -104
rect 33 -111 46 -104
rect 51 -111 59 -104
rect 64 -111 73 -104
rect 78 -111 93 -104
rect 98 -111 102 -79
rect 0 -160 7 -139
rect 141 -163 154 -3
rect 141 -188 153 -163
rect -159 -213 153 -188
<< ntransistor >>
rect -30 -25 -23 -13
rect 27 -25 34 -13
rect 88 -25 95 -13
rect -91 -82 -85 -70
rect -29 -82 -23 -70
rect 28 -81 34 -69
rect 89 -81 95 -69
<< ptransistor >>
rect -92 72 -86 84
rect -28 71 -22 83
rect 27 70 33 82
rect 88 70 94 82
rect -30 31 -23 43
rect 27 31 34 43
rect 88 31 95 43
<< polycontact >>
rect -92 39 -78 45
rect -132 -7 -126 3
rect 5 -2 11 7
rect 65 -2 71 7
rect 0 -139 7 -127
<< ndcontact >>
rect -36 -23 -32 -16
rect -20 -23 -16 -16
rect 20 -23 24 -16
rect 36 -23 40 -16
rect 82 -23 86 -16
rect 98 -23 102 -16
rect -97 -80 -93 -73
rect -82 -80 -78 -73
rect -35 -80 -31 -73
rect -21 -80 -17 -73
rect 21 -79 25 -72
rect 37 -79 41 -72
rect 82 -79 86 -72
rect 98 -79 102 -72
<< pdcontact >>
rect -97 74 -93 82
rect -82 75 -78 82
rect -36 73 -31 80
rect -21 73 -16 81
rect 20 72 24 79
rect 35 72 39 79
rect 82 72 87 79
rect 97 72 101 79
rect -36 33 -32 40
rect -20 33 -16 40
rect 20 33 24 40
rect 36 33 40 40
rect 82 33 86 40
rect 97 33 102 40
<< psubstratepcontact >>
rect -91 -111 -86 -104
rect -77 -111 -72 -104
rect -64 -111 -59 -104
rect -38 -111 -33 -104
rect -26 -111 -21 -104
rect -10 -111 -5 -104
rect 14 -111 19 -104
rect 28 -111 33 -104
rect 46 -111 51 -104
rect 59 -111 64 -104
rect 73 -111 78 -104
rect 93 -111 98 -104
<< nsubstratencontact >>
rect -100 97 -96 102
rect -90 97 -86 102
rect -81 97 -77 102
rect -38 98 -34 103
rect -30 98 -26 103
rect -15 98 -11 103
rect 15 98 19 103
rect 24 98 28 103
rect 40 98 44 103
rect 78 98 82 103
rect 87 98 91 103
rect 100 98 104 103
<< labels >>
rlabel metal1 -100 103 -99 103 5 vdd
rlabel metal1 2 -155 3 -155 1 vctrl
rlabel metal1 128 1 129 1 1 out
rlabel metal1 -96 -109 -96 -109 1 gnd
rlabel metal1 -82 7 -82 7 1 mid1
rlabel metal1 -11 2 -11 2 1 mid2
rlabel metal1 43 1 43 1 1 mid3
rlabel metal1 -35 58 -35 58 1 top1
rlabel metal1 21 58 21 58 1 top2
rlabel metal1 83 58 83 58 1 top3
rlabel metal1 -34 -50 -34 -50 1 bot1
rlabel metal1 21 -47 21 -47 1 bot2
rlabel metal1 83 -48 83 -48 1 bot3
<< end >>
